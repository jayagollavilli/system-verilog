`ifndef"ALL_INTF"
`define"ALL_INTF"
interface intf();
logic a;
logic b;
logic[6:0]c;
endinterface:intf
`endif

